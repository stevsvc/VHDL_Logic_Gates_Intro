LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY work;

ENTITY VHDL_newGates IS
	PORT
	(
		IN_1, IN_2, IN_3, IN_4, POLARITY_CNTRL: IN BIT;
		OUT_1, OUT_2, OUT_3, OUT_4: OUT BIT
	);
END VHDL_newGates;

ARCHITECTURE new_gates OF VHDL_newGates IS

BEGIN 

OUT_1 <= IN_1 NAND POLARITY_CNTRL;
OUT_2 <= IN_2 AND POLARITY_CNTRL;
OUT_3 <= IN_3 NOR POLARITY_CNTRL;
OUT_4 <= IN_4 XNOR POLARITY_CNTRL;

END new_gates;